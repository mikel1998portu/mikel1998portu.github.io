�PNG

   IHDR  @  +   &�}$   PLTE &��&   $z��C��\Hեv傅  �IDATx����o$e~��6��*Z��B!>G��(��Bp�a��\֠F�(�C�� �0?��岬4H!�J��rHX4"V��ǎm懱�ޮ����-�y�m�{����~�������]�l���	@  ��@@ �@@  ��@@ �@@  ��@ ��@@  ��@ ��@@  � ��@@  � ��@@  ��@@  ��@@  �	@  ��@@ �@@  ��@@ �@@  ��@ ��@@  ��@ ��@@  � ��@@  � ��@@  ��@@  ��@@  �	@  ��@@ �@@  ��@@ �@@  ��@ ��@@  ��@ ��@@  � ��@@  � ��@@  ��@@  ��@@  �	@  ��@@ �@@  ����6���m�Ph����xh�Bk+�AR�a��
������V�Xk��@(�i�%��L��ح���� ��1�B�����D ��Ô.��aJ�ρ��D �����u��#-�1�O�ܲ%B�����-!r�?�gK��w�aJ9� 1���� ��p�汥�ى�ᡇ�?|$D �p������9��#!�#�?L����jJ�3����Ќ>���B�nJ�ݔ.3�)] ftS�@��t���M�!0���B`F7����nJ�ݔ.B3�)] ftS�@��t���M�!��0����.�<�%S�@�.L�!�����Bho1�]B����x���'��@(�Y�Kl��(���S�!��p�P ���rf���]�S�!��p�P ��c�F �)�*��Ƕ�@8�i�|�P V9U(B�	�
³��r��@�r��@μQ60��Z{	C�@κ��73�G g\p'q�����.�T_�?n�N� �!oܙgW��h��}��o���km� ��晐�O�s @ ˚������F����,���:�ԓ+��<�
���-%2��9i�~_X}��uQ�@��y1k9��춲 ��{<zARۑw�vy�ւha��^�D϶�m���ɯ��ѯ}�۟|����Y��������������?�g3/���&� ���ן�t�o�L��O+A!��c/���Fo��/.��������$��B�;������>�����R��щ�����5v����G����{{�w'g���A3�=����iS7^�Z�qCw6ze��#��X�n�IC7�Y�n5�ǋy���=�Y���ٺ�A��Y�f�䇹}4|@ g��y_����g����F��;���@β�_o8���B�6��Y0����
K �*:Q���gD��$Z�[߰�Ȳv�.���ef�J��K��W��kw�_ �+n.YH��z,��{������]�,?�~g�ý�e��Z��GA������R����R+�T܇���	���?���/��/�ƺt�zn��k�5V�X֫��V+}��TR 6�2k���z�B��I4��PVXi}��_H���*�T�{2���#��H3§��ބ�jc��x���~�3+�F�������{�Hj������� �4�Q�B��<묱F����a[�4�ꂗ�-��j��^\�}*
�)���{�O�W�D��'�/e�7'�ͳ��ʪ: ܫ��zsѹ*
�9_�Ue�Z�T|�_p k�BE�4i�Q��'m�ޫ�Zp �Ҝ��;�j�z�ö�����8��gU �Y����5'��A�kޟY<�8�.�&�i����8�T��s%.nt] M������x�?z��� N��a%^���gCjA*��B^,�3N��YWK�Lٳ!�Z��;)�s���98�.�f�jU�5��z����a���it�4��T;��_�'�+�S/��!��ҴRS��q�:Ws@.u*��R7>�|
�a���9�U�"��BF[�nɧ�Ҵ�'�ߚ���Q�_�Pbz�ܜ2�|
�i�.^Z|�i�s���ϕ��A^�4�j��p�Wy����z���8�+��|�_t2��~x��y���y҂��/���}�>,��w�W m(����GK������7%o�g�҆sM����c�^~B�Y�*�m�W�`��r��(�ޗ�=��
����o��G'����！Yzٿ���}���� �@�q���O��eC��Q酓��x7y��8��G.������I�w���`o{��u�;�pմ�7�~�b���^����?q1�rH�@.-�/?|-�^t�o?5]x������|�?/�8���;��xnT i:����/��/��]ȃ�xTG�@x���W�i`r�!���@�	d�����x�xr��n�NK�f?�X=x����ȏ�-θī_ ��Z�|"�oϸ�H��)<嫭i�{߹���]p������W��x��Hk�)����߾]�y����[ǃF��<������z��m[3�=�����y�>��\������L�v �+�x�L�7� �@b�l�F����������;�����G_=lo��N��|������';�NS���n裯��L��	Ҧ�ٸy�U�f�GWr�����+�6����8�������+�6�߀o�����yҦ�;�(�G܍�x�@�|�K�gt&H��o�u��y�SRV����/�܎� ��j�H�!������� �30�����D q��q��� �@�BƵ߿�p�"���뿁w�e#�@����xF�D q�߆#!{F�D����iHl���sq۶D �?w��cAb�=���99�CHx��	�!�ħmrƇ��2��	�l!F��?�D<�{���@�B�D���&������F�$?�D<_�fH�CHĥL��M ��$�2�Dwl1���'��υX��^݅N��If+�3(���h��tZ~M=k��v��K�eH���+�X�"�.=^w�Ӣ�D �!�o��<�]#�@����>3u/ŹH ��TLR��b9����f5wx��!$�!յ~��rf��H뙬���t=��c<��D 	�\�f�"������A��Ї��\�8���C �\��Z��i�ǉ�āe�+ҽ�nb����v�@ g\h71���.U�z�ҽ��z��N
$�E���iB��0�����k��H�EM��kI��B�Ta�EM���L �ߴ']?�QR�3�0=������8M(�8zr�t�3%�(��']?�M3�@�S|�t��2��~N �P��`�Vg?�@Z5L�UY����$�H��q*���k�f�Β��T�&H�Sz��)^����IqJ��c�3�@z5�w|�wVc'�@�-�;>�[<�{������ʦp���$�)}�����ҳ)��K����ٔ��.�Ĝҳ.�܌.��M��[�ft��l	��q�53�@Ҵ��t�������ߙt� F��^��k�Yw���׺$�y���y+I)U��,�J��IvJ�����] ���;|�^3��Szw�� �Pm���p1�<�@�G_��������3�@�37�$]�'�:�֓�o����o��hдY�72ώ@�۩\NWS�M���c��E;
������?�.T ^l2���w#߿@ګ:tu��A,��`^u68e�/��U��fM
�� �@Ұ]u8h֬���t*��
-uv<3I°�p�M�cό@��Ru:hԨ��tk��tШ�Ig�H�1�Ë�_�{^�����A��Z�$.�bfRu�@:6���F�*��H�V*~�����XIE��L��O �X���@�+����xs@Q>N(�td��?>N(�t��Ǟ�$c/ޞe^qՇ@�W�*��#S��V}�䂦��Lͪ-�H��&��U[�!�֫-��yb��ij�Ǟ�$��j�Is��V��&$���^�Sω@R2�4B7gn�%�>(8�����I���HZ
v��)�Uڱ �H��f�ƬUZ�!HzV"-u�J;�N�!�)E����e\i�n�n���D�e�S��s�W �Y��
�b�JCtS��&"˰�ݐI���D�Wi�nʬ�@�@��W����ea'�KhY�(�@z�ciJVe��@"�qu�ȳ*���FXyp�W 鉱�_I~�������,�!�u�] �I�S�Sφ@ғ��o�Z�I2Ӑ@���kMf��@z#4n�Z����R �8�W�4�@��&Ƕ�@��l<���g
'�C$�m9k�w���ٸ�kM�H�$2;O(�4mw���W��Hd�S�Pl�����N��B$���c�R�BlkF![�t�X�@��1�
_E ��O����@�2�**@ ���uû&!_��#�w{w+�R���4����8'������y
G
2�@ �� Ҥ�����W+�{�������yg� �3g-���q�]�+��]i"�tu; g�Q��K�����N��C~3�@�&��$�qr�����CH�v�,��+M�7�^�n{��,6�,$Y�c��Rr:dޗK����M �0���K���܃�Ny��wx_3O�@�f���.Oy�VQ  ���=���G
sOЏ=��S����U�`I@�ׄ�6V����{bcuZ���q���i�#���j�i8���'6��f�F�W�<z�8�ĭ\����]�kwn����w��ֿ��.f^� �6�n�W���S��^`��@zm2���*h��bk��H���V'�Guܩ��8>�\�|�a#>�.���Sz��.ԯ������OM������o}�����{�1����`�o��] =t�g�w�������lW��7��y�M�2�a6h���޽�����M }4�	�4G=��|^J is*[ �k�&���Z�6�@��Z��@�#�)���M  �S�y|��@z������mܺM �J0��@zljB��m��@��G293\J,�l�`"ȩ�c�!`�&� �Ú�#��C��~�����ҭ����h���jfc	�����t�����kw�"�Yqyo�T�*yg?�;���:�<9����\���p�ȩ��ڻ����<޸jd�&H��ŧ�K��;�Z�Ǌ���i3룃��Fr����ﳭoo��7���YYm5~�ǵ�;���}����*wf��H���j���Zo}���1�o��:���N�H�;?�{r���]$��V�b`���V�.߱���rw��@@   ��@@   ��@@  @  ��@@  @  ��@@ �@@  ��@@ �@@  ��@ ��@@  ��@ ��@@  � ��@@  � ��@@  � ��@@  ��@@  Um��~i؃�@@  @  ��@@  @  ��@@ �@@  ��@@ �@@  ��@@ 6��@@  ��@@  ��@@   ��@@   ��@@  @  ��@@  @  ��@@ �@@  ��@@ �@@  ��@@ 6��@@  ��@@  ��@@   ��@@   ��@@  @  ��@@  @  ��@@ �@@  ��@@ �@@  ��@@ 6��@@  ��@@  ��@@   ��@@   ��@@  @  ��@@  @  h�����-y��    IEND�B`�